//
// Copyright 2009 Erik Gilling
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//

module ir(
    output reg [7:0] ir,
    input [7:0]      data,
    input 	     sync,
    input 	     rst_n);

   always @(posedge sync or negedge rst_n) begin
      if (rst_n == 1'b0) begin
	 ir = 8'h00;
      end else if (sync == 1'b1) begin
	 ir = data;
      end
   end
endmodule
      