//
// Copyright 2009 Erik Gilling
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//

`timescale 1ns/1ps

module sram (
    inout [7:0] data,
    input [10:0] 	addr,
    input 		w,
    input 		oe);

   reg [7:0] 	sram[0:2048-1];

   assign data = oe == 1'b1 ? sram[addr] : 8'hZ;

   always @(posedge w) begin
      sram[addr] <= data;
   end
endmodule
