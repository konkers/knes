`timescale 1ns / 1ps

// 6502 toplevel module.
module k6502(
    inout [7:0] d,
    inout [15:0] a,
    input reset_n,
    input ph0,
    output ph1_out,
    output ph2_out
);

wire ph1;
wire ph2;
clockgen clockgen(
    .ph0(ph0),
    .ph1(ph1),
    .ph2(ph2),
    .ph1_out(ph1_out),
    .ph2_out(ph2_out)
);

control_signals_t ctl;

control_signals control_signals(ctl);
k6502_data data_half(d, a, ph1, ph2, ctl);
    

endmodule